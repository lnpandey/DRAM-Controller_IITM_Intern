package p1

endpackage : p1
